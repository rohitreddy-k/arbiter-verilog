module arbiter();
	wire S_1,S_2,S_3;
	wire 

